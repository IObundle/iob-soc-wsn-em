//mixer 
`define LPF_ADDR_W 1

`define LPF_PD 0
`define LPF_FC 1

