//mixer 
`define MIXER_ADDR_W 2

`define MIXER_PD 0
`define MIXER_OTA 1
`define MIXER_BUFF 2

