`timescale 1ns / 1ps


///////////////////////////////////////////////////////////////////////////////
// Date: 26/09/2020
// Module: limiter.sv
// Project: WSN
// Description: emulates the limiter behaviour
//				 


module limiter(input real signal_in, output bit square_out, input limiter_pd);


   parameter offset = 0;
   
   //-------------------------------- Signal Limiting---- -------------------------------
   assign square_out = limiter_pd ? 0 : ((signal_in > offset)? 1 : 0);

   
endmodule

