//iref
`define IREF_ADDR_W 1

`define IREF_PD (`IREF_ADDR_W'd0)
`define IREF_FC (`IREF_ADDR_W'd1)

