
   pa_tb pa_tb0
     (
      .in      (pa_i),
      .out     (pa_o),
      .pd      (pa_pd),
      .mode    (pa_mode)
      );

