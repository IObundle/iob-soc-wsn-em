//pa 
`define PA_ADDR_W 1

`define PA_PD   (`PA_ADDR_W'd0)
`define PA_MODE (`PA_ADDR_W'd1)

