//pa 
`define PA_ADDR_W 1

`define PA_PD 0
`define PA_MODE 1

