`define TMP_ADDR_W 1

`define TMP_VALUE (`TMP_ADDR_W'd0)   //Read

`define ADC_RESOLUTION 10            //ADC resolution 
`define RDATA_W        32            //rdata width

`define RDATA_RVAL     32'b0         //rdata reset value  
