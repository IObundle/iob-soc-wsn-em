// ID
`define ID_ADDR_W 1

`define ID_VALUE (`ID_ADDR_W'd0)
