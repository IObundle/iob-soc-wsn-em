
   pa_tb pa_tb0
     (
      .in      (pa_io),
      .out     (pa_io),
      .pd      (pa_pd),
      .mode    (pa_mode)
      );

