//mixer 
`define MIXER_ADDR_W 2

`define MIXER_PD   (`MIXER_ADDR_W'd0)
`define MIXER_OTA  (`MIXER_ADDR_W'd1)
`define MIXER_BUFF (`MIXER_ADDR_W'd2)

