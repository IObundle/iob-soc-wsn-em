
   lna_tb lna_tb0
     (
      .lna_in      (lna_io_tb),
      .lna_out     (lna_io_tb),
      .lna_pd      (lna_pd_tb),
      .lna_mode    (lna_mode_tb)
      );

