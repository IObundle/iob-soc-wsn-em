
   iref_tb iref_tb0
     (
      .charge       (iref_charge_tb),
      .pd           (iref_pd_tb)
      );

