//lpf
`define LPF_ADDR_W 1

`define LPF_PD (`LPF_ADDR_W'd0)
`define LPF_FC (`LPF_ADDR_W'd1)

