`define LIMITER_ADDR_W 1

`define LIMITER_PD (`LIMITER_ADDR_W'd0)
