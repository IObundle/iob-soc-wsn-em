
   lpf_tb lpf_tb0
     (
      .sampling_clk (lpf_sampling_clk_tb),
      .in           (lpf_in_tb),
      .out          (lpf_out_tb),
      .fc           (lpf_fc_tb),
      .pd           (lpf_pd_tb)
      );

