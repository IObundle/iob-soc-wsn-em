//iref
`define IREF_ADDR_W 1

`define IREF_PD 0
`define IREF_FC 1

