
   pa_tb pa_tb0
     (
      .in      (pa_io_tb),
      .out     (pa_io_tb),
      .pd      (pa_pd_tb),
      .mode    (pa_mode_tb)
      );

