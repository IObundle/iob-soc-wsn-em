//lna 
`define LNA_ADDR_W 1

`define LNA_PD 0
`define LNA_MODE 1

